��Q      �sklearn.linear_model._logistic��LogisticRegression���)��}�(�penalty��l2��dual���tol�G?6��C-�C�G?�      �fit_intercept���intercept_scaling�K�class_weight�N�random_state�N�solver��lbfgs��max_iter�Kd�multi_class��auto��verbose�K �
warm_start���n_jobs�N�l1_ratio�N�feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�P1��P2��P4��P5��P6�et�b�n_features_in_�K�classes_�hhK ��h��R�(KK��h$�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�n_iter_�hhK ��h��R�(KK��h$�i4�����R�(Kh:NNNJ����J����K t�b�C   �t�b�coef_�hhK ��h��R�(KKK��h$�f8�����R�(Kh:NNNJ����J����K t�b�C(-Do@h��?T�\���?���f����"��Y�?Fֵ����?�t�b�
intercept_�hhK ��h��R�(KK��hP�C-�8�VO ��t�b�_sklearn_version��1.1.1�ub.